module cla_32_bit_adder(
            A,
            B,
            Cin,
            S_reg,
            Cout_reg,
            clk);
    input clk;
    input [31:0] A, B;
    input Cin;
    wire [7:0] C;
    wire [7:0] P, G;
    wire [31:0] S;
    reg Cout;

    reg [31:0] A_reg, B_reg;
	reg Cin_reg;
	output reg [31:0] S_reg;
	output reg Cout_reg;

    // registers
    always @ (posedge clk) begin
        A_reg <= A;
        B_reg <= B;
        Cin_reg <= Cin;
        S_reg <= S;
        Cout_reg <= C[7];
    end

    cla_32_bit_module cla (Cin_reg, P, G, C);

    cla_4_bit_adder c0 (A_reg[3:0],
                B_reg[3:0],
                Cin_reg,
                S[3:0],
                P[0],
                G[0]);

    cla_4_bit_adder c1 (A_reg[7:4],
                B_reg[7:4],
                C[0],
                S[7:4],
                P[1],
                G[1]);

    cla_4_bit_adder c2 (A_reg[11:8],
                B_reg[11:8],
                C[1],
                S[11:8],
                P[2],
                G[2]);

    cla_4_bit_adder c3 (A_reg[15:12],
                B_reg[15:12],
                C[2],
                S[15:12],
                P[3],
                G[3]);

    cla_4_bit_adder c4 (A_reg[19:16],
                B_reg[19:16],
                C[3],
                S[19:16],
                P[4],
                G[4]);

    cla_4_bit_adder c5 (A_reg[23:20],
                B_reg[23:20],
                C[4],
                S[23:20],
                P[5],
                G[5]);

    cla_4_bit_adder c6 (A_reg[27:24],
                B_reg[27:24],
                C[5],
                S[27:24],
                P[6],
                G[6]);

    cla_4_bit_adder c7 (A_reg[31:28],
                B_reg[31:28],
                C[6],
                S[31:28],
                P[7],
                G[7]);




    // always @ * begin
        // C[0] = Cin_reg;
        // C[1] <= Cin_reg & P[0] | C[0];
        // C[2] <= G[0] & P[1] | C[1];
        // C[3] <= G[1] & P[2] | C[2];
        // C[4] <= G[2] & P[3] | C[3];
        // C[5] <= G[3] & P[4] | C[4];
        // C[6] <= G[4] & P[5] | C[5];
        // C[7] <= G[5] & P[6] | C[6];
        // Cout <= G[6] & P[7] | C[7];
        // // C[1] = (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))));
        // // C[2] = (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))));
        // // C[3] = (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))));
        // // C[4] = (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))));
        // // C[5] = (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))));
        // // C[6] = (G[23] | P[23] & (G[22] | P[22] & (G[21] | P[21] & (G[20] | P[20] & (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))))))));
        // // C[7] = (G[27] | P[27] & (G[26] | P[26] & (G[25] | P[25] & (G[24] | P[24] & (G[23] | P[23] & (G[22] | P[22] & (G[21] | P[21] & (G[20] | P[20] & (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))))))))))));
        // // Cout = (G[31] | P[31] & (G[30] | P[30] & (G[29] | P[29] & (G[28] | P[28] & (G[27] | P[27] & (G[26] | P[26] & (G[25] | P[25] & (G[24] | P[24] & (G[23] | P[23] & (G[22] | P[22] & (G[21] | P[21] & (G[20] | P[20] & (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))))))))))))))));
    // end


    // generate
    //     genvar j;
    //     for (j = 0; j < 32; j = j + 1) begin : jate
    //         assign C[j + 1] = G[j] | P[j] & C[j];
    //     end
    // endgenerate

    // assign

        // C[0] <= Cin_reg;
        // C[1] <= Cin_reg & P[0] | G[0];
        // C[2] <= G[0] & P[1] | G[1];
        // C[3] <= G[1] & P[2] | G[2];
        // C[4] <= G[2] & P[3] | G[3];
        // C[5] <= G[3] & P[4] | G[4];
        // C[6] <= G[4] & P[5] | G[5];
        // C[7] <= G[5] & P[6] | G[6];
        // Cout <= G[6] & P[7] | G[7];
        // C[1] <= (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))));
        // C[2] <= (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))));
        // C[3] <= (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))));
        // C[4] <= (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))));
        // C[5] <= (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))));
        // C[6] <= (G[23] | P[23] & (G[22] | P[22] & (G[21] | P[21] & (G[20] | P[20] & (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))))))));
        // C[7] <= (G[27] | P[27] & (G[26] | P[26] & (G[25] | P[25] & (G[24] | P[24] & (G[23] | P[23] & (G[22] | P[22] & (G[21] | P[21] & (G[20] | P[20] & (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))))))))))));
        // Cout <= (G[31] | P[31] & (G[30] | P[30] & (G[29] | P[29] & (G[28] | P[28] & (G[27] | P[27] & (G[26] | P[26] & (G[25] | P[25] & (G[24] | P[24] & (G[23] | P[23] & (G[22] | P[22] & (G[21] | P[21] & (G[20] | P[20] & (G[19] | P[19] & (G[18] | P[18] & (G[17] | P[17] & (G[16] | P[16] & (G[15] | P[15] & (G[14] | P[14] & (G[13] | P[13] & (G[12] | P[12] & (G[11] | P[11] & (G[10] | P[10] & (G[9] | P[9] & (G[8] | P[8] & (G[7] | P[7] & (G[6] | P[6] & (G[5] | P[5] & (G[4] | P[4] & (G[3] | P[3] & (G[2] | P[2] & (G[1] | P[1] & (G[0] | P[0] & Cin_reg))))))))))))))))))))))))))))))));




    // cla_4_bit c0 (A_reg[3:0],
    //             B_reg[3:0],
    //             C[0],
    //             S[3:0],
    //             P[3:0],
    //             G[3:0],
    //             C[4]);
    //
    // cla_4_bit c1 (A_reg[7:4],
    //             B_reg[7:4],
    //             C[4],
    //             S[7:4],
    //             P[7:4],
    //             G[7:4],
    //             C[8]);
    //
    // cla_4_bit c2 (A_reg[11:8],
    //             B_reg[11:8],
    //             C[8],
    //             S[11:8],
    //             P[11:8],
    //             G[11:8],
    //             C[12]);
    //
    // cla_4_bit c3 (A_reg[15:12],
    //             B_reg[15:12],
    //             C[12],
    //             S[15:12],
    //             P[15:12],
    //             G[15:12],
    //             C[16]);
    //
    // cla_4_bit c4 (A_reg[19:16],
    //             B_reg[19:16],
    //             C[16],
    //             S[19:16],
    //             P[19:16],
    //             G[19:16],
    //             C[20]);
    //
    // cla_4_bit c5 (A_reg[23:20],
    //             B_reg[23:20],
    //             C[20],
    //             S[23:20],
    //             P[23:20],
    //             G[23:20],
    //             C[24]);
    //
    // cla_4_bit c6 (A_reg[27:24],
    //             B_reg[27:24],
    //             C[24],
    //             S[27:24],
    //             P[27:24],
    //             G[27:24],
    //             C[28]);
    //
    // cla_4_bit c7 (A_reg[31:28],
    //             B_reg[31:28],
    //             C[28],
    //             S[31:28],
    //             P[31:28],
    //             G[31:28],
    //             C[32]);


    // integer j;
    // always @ (*) begin
    //     for (j = 0; j < 32; j = j + 1) begin : jate
    //         C[j + 1] = G[j] | P[j] & C[j];
    //         end
    // end
    //
    // generate
    //     genvar i;
    //     for (i = 0; i < 8; i = i + 1) begin : nate
    //         cla_4_bit c (A_reg[(i + 1) * 4 - 1:i * 4],
    //                     B_reg[(i + 1) * 4 - 1:i * 4],
    //                     C[(i + 1) * 4 - 1:i * 4],
    //                     S[(i + 1) * 4 - 1:i * 4],
    //                     P[(i + 1) * 4 - 1:i * 4],
    //                     G[(i + 1) * 4 - 1:i * 4]);
    //         end
    // endgenerate

endmodule
